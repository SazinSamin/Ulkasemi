`timescale 1ns/1ps

module counter(
  input [15:0] data_in,
  input load,
  input enable,
  input up_down,
  input clk,
  input reset,
  output wire [15:0] data_out
);






endmodule