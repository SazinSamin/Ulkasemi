package counter_tb_package;
  `include "counter_stimulus.sv";
  `include "counter_driver.sv";
  `include "counter_monitor.sv";
  `include "counter_agent.sv";
  `include "counter_scoreboard.sv";  
  `include "counter_environment.sv";
  `include "counter_test.sv"
endpackage 