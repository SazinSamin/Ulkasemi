class counter_scoreboard;

  function new();
    $display("%0t Counter_Scoreboard Created", $time);
  endfunction : new


endclass