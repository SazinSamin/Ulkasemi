module counter(
  input [15:0] data_in,
  input load,
  input enable,
  input up_down,
  input clk,
  input reset,
  output [15:0] data_out
);
endmodule