class counter_driver;

  function new(virtual counter_interface count_vif);
    $display("driver class created successfully");
  endfunction

endclass