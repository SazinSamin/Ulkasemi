class counter_scoreboard;
  
  function new();
    $display("scoreboard class created successfully");

  endfunction
endclass