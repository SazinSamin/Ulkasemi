class counter_monitor;

  function new();
    $display("monitor class created successfully");
  endfunction
  
endclass